`default_nettype none
`timescale 1ns/1ns

// ARITHMETIC-LOGIC UNIT
// > Executes computations on register values
// > In this minimal implementation, the ALU supports the 4 basic arithmetic operations
// > Each thread in each core has it's own ALU
// > ADD, SUB, MUL, DIV instructions are all executed here
module alu (
    input  wire         clk,
    input  wire         reset,
    input  wire         enable, // If current block has less threads then block size, some ALUs will be inactive

    input  reg  [2:0]   core_state,

    input  reg  [1:0]   decoded_alu_arithmetic_mux,
    input  reg          decoded_alu_output_mux,

    input  reg  signed [7:0]   rs,
    input  reg  signed [7:0]   rt,
    output reg  [7:0]          alu_out
);
    localparam ADD = 2'b00,
               SUB = 2'b01,
               MUL = 2'b10,
               DIV = 2'b11;

    always @(posedge clk) begin 
        if (reset) begin 
            alu_out <= 8'b0;
        end else if (enable) begin
            // Calculate alu_out when core_state = EXECUTE
            if (core_state == 3'b101) begin 
                if (decoded_alu_output_mux == 1) begin 
                    // Set values to compare with NZP register in alu_out[2:0]
                    //mofify to signed calculation
                    alu_out <= {5'b0, ($signed(rs) - $signed(rt) > 0), ($signed(rs) - $signed(rt) == 0), ($signed(rs) - $signed(rt) < 0)};
                end else begin 
                    // Execute the specified arithmetic instruction
                    case (decoded_alu_arithmetic_mux)
                        ADD: begin 
                            alu_out <= rs + rt;
                        end
                        SUB: begin 
                            alu_out <= rs - rt;
                        end
                        MUL: begin 
                            alu_out <= rs * rt;
                        end
                        DIV: begin 
                            alu_out <= rs / rt;
                        end
                    endcase
                end
            end
        end
    end
endmodule
